module seven_segment(in0,in1,op_code,enable,a,b,c,d,e,f,g);
parameter N = 4;
input [N-1:0]in0;
input [N-1:0]in1;
input [N-3:0]op_code;
input enable;
output reg a ;
output reg b ;
output reg c ;
output reg d ;
output reg e ;
output reg f ;
output reg g ;
always @(*) begin
    if(enable==1'b1)begin
        case(op_code)
        2'b00:case (in0+in1)
          4'b0000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end   
          4'b0001:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end     
          4'b0010:begin
             a=1'b1;
             b=1'b1;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end 
          4'b0011:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b0;
             g=1'b1;
             end      
          4'b0100:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b0101:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end 
          4'b0110:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b0111:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end
          4'b1000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1001:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b1010:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1011:begin
             a=1'b0;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1100:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end
          4'b1101:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end 
          4'b1110:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1111:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          endcase              
        2'b01:case (in0|in1)
          4'b0000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end   
          4'b0001:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end     
          4'b0010:begin
             a=1'b1;
             b=1'b1;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end 
          4'b0011:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b0;
             g=1'b1;
             end      
          4'b0100:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b0101:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end 
          4'b0110:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b0111:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end
          4'b1000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1001:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b1010:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1011:begin
             a=1'b0;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1100:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end
          4'b1101:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end
          4'b1110:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1111:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
           endcase
        2'b10:case (in0-in1)
          4'b0000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end   
          4'b0001:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end     
          4'b0010:begin
             a=1'b1;
             b=1'b1;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end 
          4'b0011:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b0;
             g=1'b1;
             end      
          4'b0100:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b0101:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end 
          4'b0110:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b0111:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end
          4'b1000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1001:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b1010:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1011:begin
             a=1'b0;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1100:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end
          4'b1101:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end
          4'b1110:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1111:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          endcase
        2'b11:case (in0^in1)
          4'b0000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end   
          4'b0001:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end     
          4'b0010:begin
             a=1'b1;
             b=1'b1;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end 
          4'b0011:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b0;
             g=1'b1;
             end      
          4'b0100:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b0101:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end 
          4'b0110:begin
             a=1'b1;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b0111:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b0;
             f=1'b0;
             g=1'b0;
             end
          4'b1000:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1001:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b0;
             f=1'b1;
             g=1'b1;
             end
          4'b1010:begin
             a=1'b1;
             b=1'b1;
             c=1'b1;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1011:begin
             a=1'b0;
             b=1'b0;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1100:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b0;
             end
          4'b1101:begin
             a=1'b0;
             b=1'b1;
             c=1'b1;
             d=1'b1;
             e=1'b1;
             f=1'b0;
             g=1'b1;
             end
          4'b1110:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b1;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end
          4'b1111:begin
             a=1'b1;
             b=1'b0;
             c=1'b0;
             d=1'b0;
             e=1'b1;
             f=1'b1;
             g=1'b1;
             end                                                                   
          endcase
        endcase
        end
     else if(enable==1'b0) begin
            
        end
end
endmodule
